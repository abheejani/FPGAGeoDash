module Rand(input Clk, input Reset, input str,
				output [10:0] randNum1,randNum2,randNum3
);

		
endmodule 